library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity WB_Register is 
    Port ( Clk, Rst, WE, Din_1, Din_2 : in  std_logic;
           Dout_1, Dout_2 			  : out std_logic
	);
end WB_Register;

architecture Behavioral of WB_Register is

begin


end Behavioral;

